`timescale 1ns/1ns


`define X_LENGTH 32

`define REGISTER_WIDTH 5
`define REGISTER_COUNT 32

`define MEMORY_WIDTH 32
`define MEMORY_DEPTH 5
`define MEMORY_COUNT 32

// `define DECODE_INFO_WIDTH (10 + 9 + 6 + 2 + 2 + 3 + 5 + 8 + 2)
